// No work done here yet, just a placeholder for the future.